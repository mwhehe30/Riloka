<svg width="88" height="88" viewBox="0 0 88 88" fill="none" xmlns="http://www.w3.org/2000/svg">
  <defs>
    <linearGradient id="grad" x1="0" y1="0" x2="88" y2="88" gradientUnits="userSpaceOnUse">
      <stop stop-color="#6366F1"/>
      <stop offset="1" stop-color="#06B6D4"/>
    </linearGradient>
    <linearGradient id="grad2" x1="44" y1="20" x2="44" y2="70" gradientUnits="userSpaceOnUse">
      <stop stop-color="#FB7185"/>
      <stop offset="1" stop-color="#F9A8D4"/>
    </linearGradient>
  </defs>
  <circle cx="44" cy="44" r="40" fill="url(#grad)" opacity="0.1"/>
  <path d="M44 18C31 18 20 29 20 42C20 51 26 59 33 65L44 76L55 65C62 59 68 51 68 42C68 29 57 18 44 18ZM44 46C40.69 46 38 43.31 38 40C38 36.69 40.69 34 44 34C47.31 34 50 36.69 50 40C50 43.31 47.31 46 44 46Z" fill="url(#grad)"/>
  <circle cx="44" cy="40" r="5" fill="url(#grad2)"/>
</svg>
